    Mac OS X            	   2  �     �                                    ATTR     �   �  �                  �  �  #com.apple.fileutil.PlaceholderData   DENO      �                     `                7d6b03d2adf04fc0b2a7227ce46c6525        7d6b03d2adf04fc0b2a7227ce46c6525        b7c075b82d074e23949a0b803d2bb1a4       423ea328676e43ccb769dfb6a5e7ea8d        25ec87dd70c745fcb3a5603859fcf0bc        c849699375d54c8e84bca7a577bc1431        c475ffdd-e381-471e-b27d-50cda663f7a0 �U@�-�YR�9�!l<b��9�   @�-�YR�9�!l<b��9�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          This resource fork intentionally left blank                                                                                                                                                                                                                            ��